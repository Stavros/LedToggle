-- ledtoggle_tb.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ledtoggle_tb is
end entity ledtoggle_tb;

architecture rtl of ledtoggle_tb is
	component ledtoggle is
		port (
			clk_clk        : in  std_logic                    := 'X';             -- clk
			led_pin_export : out std_logic_vector(7 downto 0);                    -- export
			reset_reset_n  : in  std_logic                    := 'X';             -- reset_n
			sw_pin_export  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- export
			uart_pins_rxd  : in  std_logic                    := 'X';             -- rxd
			uart_pins_txd  : out std_logic                                        -- txd
		);
	end component ledtoggle;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_conduit_bfm is
		port (
			sig_export : in std_logic_vector(7 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm_0002 is
		port (
			sig_export : out std_logic_vector(7 downto 0)   -- export
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			sig_rxd : out std_logic_vector(0 downto 0);                    -- rxd
			sig_txd : in  std_logic_vector(0 downto 0) := (others => 'X')  -- txd
		);
	end component altera_conduit_bfm_0003;

	signal ledtoggle_inst_clk_bfm_clk_clk           : std_logic;                    -- ledtoggle_inst_clk_bfm:clk -> [ledtoggle_inst:clk_clk, ledtoggle_inst_reset_bfm:clk]
	signal ledtoggle_inst_led_pin_export            : std_logic_vector(7 downto 0); -- ledtoggle_inst:led_pin_export -> ledtoggle_inst_led_pin_bfm:sig_export
	signal ledtoggle_inst_sw_pin_bfm_conduit_export : std_logic_vector(7 downto 0); -- ledtoggle_inst_sw_pin_bfm:sig_export -> ledtoggle_inst:sw_pin_export
	signal ledtoggle_inst_uart_pins_txd             : std_logic;                    -- ledtoggle_inst:uart_pins_txd -> ledtoggle_inst_uart_pins_bfm:sig_txd
	signal ledtoggle_inst_uart_pins_bfm_conduit_rxd : std_logic_vector(0 downto 0); -- ledtoggle_inst_uart_pins_bfm:sig_rxd -> ledtoggle_inst:uart_pins_rxd
	signal ledtoggle_inst_reset_bfm_reset_reset     : std_logic;                    -- ledtoggle_inst_reset_bfm:reset -> ledtoggle_inst:reset_reset_n

begin

	ledtoggle_inst : component ledtoggle
		port map (
			clk_clk        => ledtoggle_inst_clk_bfm_clk_clk,              --       clk.clk
			led_pin_export => ledtoggle_inst_led_pin_export,               --   led_pin.export
			reset_reset_n  => ledtoggle_inst_reset_bfm_reset_reset,        --     reset.reset_n
			sw_pin_export  => ledtoggle_inst_sw_pin_bfm_conduit_export,    --    sw_pin.export
			uart_pins_rxd  => ledtoggle_inst_uart_pins_bfm_conduit_rxd(0), -- uart_pins.rxd
			uart_pins_txd  => ledtoggle_inst_uart_pins_txd                 --          .txd
		);

	ledtoggle_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => ledtoggle_inst_clk_bfm_clk_clk  -- clk.clk
		);

	ledtoggle_inst_led_pin_bfm : component altera_conduit_bfm
		port map (
			sig_export => ledtoggle_inst_led_pin_export  -- conduit.export
		);

	ledtoggle_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => ledtoggle_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => ledtoggle_inst_clk_bfm_clk_clk        --   clk.clk
		);

	ledtoggle_inst_sw_pin_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export => ledtoggle_inst_sw_pin_bfm_conduit_export  -- conduit.export
		);

	ledtoggle_inst_uart_pins_bfm : component altera_conduit_bfm_0003
		port map (
			sig_rxd    => ledtoggle_inst_uart_pins_bfm_conduit_rxd, -- conduit.rxd
			sig_txd(0) => ledtoggle_inst_uart_pins_txd              --        .txd
		);

end architecture rtl; -- of ledtoggle_tb
